//defines the address bus width.
`define ADDR_BUS_WIDTH 32

//defines the data bus width in terms of bytes.
`define DATA_BUS_BYTES 4

//defines the maximum write outstanding transaction capability
`define MAXWBURSTS 15

//defines the maximum read outstanding transaction capability
`define MAXRBURSTS 15
